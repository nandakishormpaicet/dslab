$date
	Sun May 23 19:23:40 2021
$end
$version
	Icarus Verilog
$end
$timescale
	1s
$end
$scope module gtob_test $end
$var wire 4 ! b [3:0] $end
$var reg 4 " g [3:0] $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
b0 "
b0 !
$end
#1
b1 !
b1 "
#2
b11 !
b10 "
#3
b10 !
b11 "
#4
b111 !
b100 "
#5
b110 !
b101 "
#6
b100 !
b110 "
#7
b101 !
b111 "
#8
b1111 !
b1000 "
#9
b1110 !
b1001 "
#10
b1100 !
b1010 "
#11
b1101 !
b1011 "
#12
b1000 !
b1100 "
#13
b1001 !
b1101 "
#14
b1011 !
b1110 "
#15
b1010 !
b1111 "
#16
